module test;

  initial begin
    $display("Hello, World!");
    $finish;  // Ends the simulation
  end

endmodule
